/* 
 * AXI stream multiplier block taking 128-bit input data and 8-bit beamforming weight to apply to data
*/
module axis_adder
  #(
    parameter SDATA_WIDTH = 128,
    parameter SSAMPLE_WIDTH = 16,
    parameter WEIGHT_WIDTH = 8,
    parameter MSAMPLE_WIDTH = 16,   // SSAMPLE_WIDTH + WEIGHT_WIDTH
    parameter MDATA_WIDTH = 128     // MSAMPLE_WIDTH * SAMPLES
   ) 
    (
/*======================================BEGIN INPUTS=======================================*/
    input wire clock,
    input wire resetn,

    // this will be the multiplication factor for all 16 samples in its channel, should be <1
    input [WEIGHT_WIDTH-1:0] bWeight00_real,
    input [WEIGHT_WIDTH-1:0] bWeight00_imag,
    input [WEIGHT_WIDTH-1:0] bWeight01_real,
    input [WEIGHT_WIDTH-1:0] bWeight01_imag,
    input [WEIGHT_WIDTH-1:0] bWeight20_real,
    input [WEIGHT_WIDTH-1:0] bWeight20_imag,
    input [WEIGHT_WIDTH-1:0] bWeight21_real,
    input [WEIGHT_WIDTH-1:0] bWeight21_imag,
    
    /* all axis prefixed variables should be inferred per UG994 because of the 
     * use of the AXI standard naming convention */
    /*-------------------------Channel00 Input Real & Imag-------------------------*/
    input wire s00_axis_real_tvalid,
    output reg s00_axis_real_tready,
    input wire [SDATA_WIDTH-1:0] s00_axis_real_tdata, // 8 16-bit samples
    input wire s00_axis_real_tlast,

    input wire s00_axis_imag_tvalid,
    output reg s00_axis_imag_tready,
    input wire [SDATA_WIDTH-1:0] s00_axis_imag_tdata, // 8 16-bit samples
    input wire s00_axis_imag_tlast,
    /*-------------------------Channel01 Input Real & Imag-------------------------*/
    input wire s01_axis_real_tvalid,
    output reg s01_axis_real_tready,
    input wire [SDATA_WIDTH-1:0] s01_axis_real_tdata, // 8 16-bit samples
    input wire s01_axis_real_tlast,

    input wire s01_axis_imag_tvalid,
    output reg s01_axis_imag_tready,
    input wire [SDATA_WIDTH-1:0] s01_axis_imag_tdata, // 16 8-bit samples
    input wire s01_axis_imag_tlast,
    /*-------------------------Channel20 Input Real & Imag-------------------------*/
    input wire s20_axis_real_tvalid,
    output reg s20_axis_real_tready,
    input wire [SDATA_WIDTH-1:0] s20_axis_real_tdata, // 16 8-bit samples
    input wire s20_axis_real_tlast,

    input wire s20_axis_imag_tvalid,
    output reg s20_axis_imag_tready,
    input wire [SDATA_WIDTH-1:0] s20_axis_imag_tdata, // 16 8-bit samples
    input wire s20_axis_imag_tlast,
    /*-------------------------Channel21 Input Real & Imag-------------------------*/
    input wire s21_axis_real_tvalid,
    output reg s21_axis_real_tready,
    input wire [SDATA_WIDTH-1:0] s21_axis_real_tdata, // 16 8-bit samples
    input wire s21_axis_real_tlast,

    input wire s21_axis_imag_tvalid,
    output reg s21_axis_imag_tready,
    input wire [SDATA_WIDTH-1:0] s21_axis_imag_tdata, // 16 8-bit samples
    input wire s21_axis_imag_tlast,
    /*-------------------------Channel21 Input Real & Imag-------------------------*/
/*=======================================END INPUTS=======================================*/

/*=====================================BEGIN OUTPUTS======================================*/
    /*-------------------------Channel00 Output Real & Imag-------------------------*/
    output reg [MDATA_WIDTH-1:0] m00_axis_real_s2mm_tdata,
    output reg [(SDATA_WIDTH/8)-1:0] m00_axis_real_s2mm_tkeep,
    output reg m00_axis_real_s2mm_tlast,
    input wire m00_axis_real_s2mm_tready,
    output reg m00_axis_real_s2mm_tvalid,

    output reg [MDATA_WIDTH-1:0] m00_axis_imag_s2mm_tdata,
    output reg [(SDATA_WIDTH/8)-1:0] m00_axis_imag_s2mm_tkeep,
    output reg m00_axis_imag_s2mm_tlast,
    input wire m00_axis_imag_s2mm_tready,
    output reg m00_axis_imag_s2mm_tvalid,
    /*-------------------------Channel01 Output Real & Imag-------------------------*/
    output reg [MDATA_WIDTH-1:0] m01_axis_real_s2mm_tdata,
    output reg [(SDATA_WIDTH/8)-1:0] m01_axis_real_s2mm_tkeep,
    output reg m01_axis_real_s2mm_tlast,
    input wire m01_axis_real_s2mm_tready,
    output reg m01_axis_real_s2mm_tvalid,

    output reg [MDATA_WIDTH-1:0] m01_axis_imag_s2mm_tdata,
    output reg [(SDATA_WIDTH/8)-1:0] m01_axis_imag_s2mm_tkeep,
    output reg m01_axis_imag_s2mm_tlast,
    input wire m01_axis_imag_s2mm_tready,
    output reg m01_axis_imag_s2mm_tvalid,
    /*-------------------------Channel20 Output Real & Imag-------------------------*/
    output reg [MDATA_WIDTH-1:0] m20_axis_real_s2mm_tdata,
    output reg [(SDATA_WIDTH/8)-1:0] m20_axis_real_s2mm_tkeep,
    output reg m20_axis_real_s2mm_tlast,
    input wire m20_axis_real_s2mm_tready,
    output reg m20_axis_real_s2mm_tvalid,

    output reg [MDATA_WIDTH-1:0] m20_axis_imag_s2mm_tdata,
    output reg [(SDATA_WIDTH/8)-1:0] m20_axis_imag_s2mm_tkeep,
    output reg m20_axis_imag_s2mm_tlast,
    input wire m20_axis_imag_s2mm_tready,
    output reg m20_axis_imag_s2mm_tvalid,
    /*-------------------------Channel21 Output Real & Imag-------------------------*/
    output reg [MDATA_WIDTH-1:0] m21_axis_real_s2mm_tdata,
    output reg [(SDATA_WIDTH/8)-1:0] m21_axis_real_s2mm_tkeep,
    output reg m21_axis_real_s2mm_tlast,
    input wire m21_axis_real_s2mm_tready,
    output reg m21_axis_real_s2mm_tvalid,

    output reg [MDATA_WIDTH-1:0] m21_axis_imag_s2mm_tdata,
    output reg [(SDATA_WIDTH/8)-1:0] m21_axis_imag_s2mm_tkeep,
    output reg m21_axis_imag_s2mm_tlast,
    input wire m21_axis_imag_s2mm_tready,
    output reg m21_axis_imag_s2mm_tvalid
/*======================================END OUTPUTS=======================================*/
    );

    integer samples = SDATA_WIDTH/SSAMPLE_WIDTH;

    integer i;

    // we need bit overflow for the following 2's complement arithmetic:
    //       reg[SSAMPLE_WIDTH] * reg[WEIGHT_WIDTH] + reg2[SSAMPLE_WIDTH] * reg2[WEIGHT_WIDTH] => 
    //          we need dataBuffer of size SSAMPLE_WIDTH+WEIGHT_WIDTH+1
    // reg [SSAMPLE_WIDTH+WEIGHT_WIDTH+1-1:0]dataBuffer; // with SSAMPLE_WIDTH=16 and WEIGHT_WIDTH=8, dataBuffer needs 25 bits
    reg [SSAMPLE_WIDTH+WEIGHT_WIDTH:0]dataBuffer00_re;  reg [SSAMPLE_WIDTH+WEIGHT_WIDTH:0]dataBuffer00_im;
    reg [SSAMPLE_WIDTH+WEIGHT_WIDTH:0]dataBuffer01_re;  reg [SSAMPLE_WIDTH+WEIGHT_WIDTH:0]dataBuffer01_im;
    reg [SSAMPLE_WIDTH+WEIGHT_WIDTH:0]dataBuffer20_re;  reg [SSAMPLE_WIDTH+WEIGHT_WIDTH:0]dataBuffer20_im;
    reg [SSAMPLE_WIDTH+WEIGHT_WIDTH:0]dataBuffer21_re;  reg [SSAMPLE_WIDTH+WEIGHT_WIDTH:0]dataBuffer21_im;

    // reg [SSAMPLE_WIDTH+3-1:0]dataBuffer_Sum;
    reg [SSAMPLE_WIDTH+2:0]dataBuffer_SumRe;
    reg [SSAMPLE_WIDTH+2:0]dataBuffer_SumIm;

    // pipelining for weights to help pass timing
    reg [7:0] bw00_re = 8'd0; reg [7:0] bw00_im = 8'd0;
    reg [7:0] bw01_re = 8'd0; reg [7:0] bw01_im = 8'd0;
    reg [7:0] bw20_re = 8'd0; reg [7:0] bw20_im = 8'd0;
    reg [7:0] bw21_re = 8'd0; reg [7:0] bw21_im = 8'd0;
    
    
    always @(posedge clock) begin
        //~resetn
        if (resetn == 1'b0) begin
            // data out, valid, tread, and tlast should all be 0
            m00_axis_real_s2mm_tdata = 1'b0;   m00_axis_imag_s2mm_tdata = 1'b0;
            m00_axis_real_s2mm_tvalid = 1'b0;  m00_axis_imag_s2mm_tvalid = 1'b0;
            s00_axis_real_tready = 1'b0;       s00_axis_imag_tready = 1'b0;
            m00_axis_real_s2mm_tlast = 1'b0;   m00_axis_imag_s2mm_tlast = 1'b0;

            m01_axis_real_s2mm_tdata = 1'b0;   m01_axis_imag_s2mm_tdata = 1'b0;
            m01_axis_real_s2mm_tvalid = 1'b0;  m01_axis_imag_s2mm_tvalid = 1'b0;
            s01_axis_real_tready = 1'b0;       s01_axis_imag_tready = 1'b0;
            m01_axis_real_s2mm_tlast = 1'b0;   m01_axis_imag_s2mm_tlast = 1'b0;

            m20_axis_real_s2mm_tdata = 1'b0;   m20_axis_imag_s2mm_tdata = 1'b0;
            m20_axis_real_s2mm_tvalid = 1'b0;  m20_axis_imag_s2mm_tvalid = 1'b0;
            s20_axis_real_tready = 1'b0;       s20_axis_imag_tready = 1'b0;
            m20_axis_real_s2mm_tlast = 1'b0;   m20_axis_imag_s2mm_tlast = 1'b0;

            m21_axis_real_s2mm_tdata = 1'b0;   m21_axis_imag_s2mm_tdata = 1'b0;
            m21_axis_real_s2mm_tvalid = 1'b0;  m21_axis_imag_s2mm_tvalid = 1'b0;
            s21_axis_real_tready = 1'b0;       s21_axis_imag_tready = 1'b0;
            m21_axis_real_s2mm_tlast = 1'b0;   m21_axis_imag_s2mm_tlast = 1'b0;
        end
        else begin

            m00_axis_real_s2mm_tlast <= s00_axis_real_tlast;    m00_axis_imag_s2mm_tlast <= s00_axis_imag_tlast;
            m01_axis_real_s2mm_tlast <= s01_axis_real_tlast;    m01_axis_imag_s2mm_tlast <= s01_axis_imag_tlast;
            m20_axis_real_s2mm_tlast <= s20_axis_real_tlast;    m20_axis_imag_s2mm_tlast <= s20_axis_imag_tlast;
            m21_axis_real_s2mm_tlast <= s21_axis_real_tlast;    m21_axis_imag_s2mm_tlast <= s21_axis_imag_tlast;

            // setting beamforming weight registers for pipelining
            bw00_re <= bWeight00_real; bw00_im <= bWeight00_imag;
            bw01_re <= bWeight01_real; bw01_im <= bWeight01_imag;
            bw20_re <= bWeight20_real; bw20_im <= bWeight20_imag;
            bw21_re <= bWeight21_real; bw21_im <= bWeight21_imag;

            /*------------------------CHANNEL 00 READY/VALID------------------------*/
            if (m00_axis_real_s2mm_tready && s00_axis_real_tvalid && m00_axis_imag_s2mm_tready && s00_axis_imag_tvalid) begin
                s00_axis_real_tready = 1'b1;       s00_axis_imag_tready = 1'b1;
                // tkeep and tvalid are now high (tkeep = 16'hffff, tvalid = 1'b1)
                m00_axis_real_s2mm_tkeep <= 16'hffff;   m00_axis_imag_s2mm_tkeep <= 16'hffff;
                m00_axis_real_s2mm_tvalid <= 1'b1;      m00_axis_imag_s2mm_tvalid <= 1'b1;

                // this for loop multiplies every eight bits by bWeights (it'll loop 16 times- 1 time per sample in tdata)
                for(i=0; i<samples; i = i+1) begin
                    // this can be a non-blocking assignment because there is a blocking assignment in the incrementing of i
                    // multiply by appropriate weight, accounting for complex/real parts of weight
                    dataBuffer00_re <= bw00_re*s00_axis_real_tdata[i*SSAMPLE_WIDTH +: SSAMPLE_WIDTH]
                        + bw00_im*s00_axis_imag_tdata[i*SSAMPLE_WIDTH +: SSAMPLE_WIDTH]; 
                    // rounding real data using bit 8
                    if (dataBuffer00_re[WEIGHT_WIDTH] == 1'b0) begin
                        m00_axis_real_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= dataBuffer00_re[SSAMPLE_WIDTH+WEIGHT_WIDTH -: SSAMPLE_WIDTH];
                    end
                    else begin // if (dataBuffer[WEIGHT_WIDTH] == 1'b1) 
                        case (dataBuffer00_re[SSAMPLE_WIDTH+WEIGHT_WIDTH -: SSAMPLE_WIDTH])
                            16'hFFFF: m00_axis_real_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= 16'hFFFF;
                            16'hEFFF: m00_axis_real_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= 16'hEFFF;
                            default:  m00_axis_real_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= dataBuffer00_re[SSAMPLE_WIDTH+WEIGHT_WIDTH -: SSAMPLE_WIDTH] + 1'b1;
                        endcase
                    end

                    dataBuffer00_im <= bw00_im*s00_axis_real_tdata[i*SSAMPLE_WIDTH +: SSAMPLE_WIDTH]
                        + bw00_re*s00_axis_imag_tdata[i*SSAMPLE_WIDTH +: SSAMPLE_WIDTH];
                    // rounding imaginary data using bit 8
                    if (dataBuffer00_im[WEIGHT_WIDTH] == 1'b0) begin
                        m00_axis_imag_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= dataBuffer00_im[SSAMPLE_WIDTH+WEIGHT_WIDTH -: SSAMPLE_WIDTH];
                    end
                    else begin // if (dataBuffer[WEIGHT_WIDTH] == 1'b1) 
                        case (dataBuffer00_im[SSAMPLE_WIDTH+WEIGHT_WIDTH -: SSAMPLE_WIDTH])
                            16'hFFFF: m00_axis_imag_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= 16'hFFFF;
                            16'hEFFF: m00_axis_imag_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= 16'hEFFF;
                            default:  m00_axis_imag_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= dataBuffer00_im[SSAMPLE_WIDTH+WEIGHT_WIDTH -: SSAMPLE_WIDTH] + 1'b1;
                        endcase
                    end
                end
            end
            /*----------------------CHANNEL 00 NOT READY/VALID----------------------*/
            else begin 
                s00_axis_real_tready = 1'b0;       s00_axis_imag_tready = 1'b0;

                // invalid data, so output data is set to static value of 0
                m00_axis_real_s2mm_tdata <= 128'b0;
                m00_axis_imag_s2mm_tdata <= 128'b0;

                // output valid and output tkeep should be low
                m00_axis_real_s2mm_tvalid <= 1'b0; m00_axis_imag_s2mm_tvalid <= 1'b0;
                m00_axis_real_s2mm_tkeep <= 1'b0;  m00_axis_imag_s2mm_tkeep <= 1'b0;
            end
            /*------------------------CHANNEL 01 READY/VALID------------------------*/
            if (m01_axis_real_s2mm_tready && s01_axis_real_tvalid && m01_axis_imag_s2mm_tready && s01_axis_imag_tvalid) begin
                s01_axis_real_tready = 1'b1;       s01_axis_imag_tready = 1'b1;
                // tkeep and tvalid are now high (tkeep = 16'hffff, tvalid = 1'b1)
                m01_axis_real_s2mm_tkeep <= 16'hffff;   m01_axis_imag_s2mm_tkeep <= 16'hffff;
                m01_axis_real_s2mm_tvalid <= 1'b1;      m01_axis_imag_s2mm_tvalid <= 1'b1;

                // this for loop multiplies every eight bits by bWeights (it'll loop 16 times- 1 time per sample in tdata)
                for(i=0; i<samples; i = i+1) begin
                    // this can be a non-blocking assignment because there is a blocking assignment in the incrementing of i
                    // multiply by appropriate weight, accounting for complex/real parts of weight
                    dataBuffer01_re <= bw01_re*s01_axis_real_tdata[i*SSAMPLE_WIDTH +: SSAMPLE_WIDTH]
                        + bw01_im*s01_axis_imag_tdata[i*SSAMPLE_WIDTH +: SSAMPLE_WIDTH]; 
                    // rounding real data using bit 8
                    if (dataBuffer01_re[WEIGHT_WIDTH] == 1'b0) begin
                        m01_axis_real_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= dataBuffer01_re[SSAMPLE_WIDTH+WEIGHT_WIDTH -: SSAMPLE_WIDTH];
                    end
                    else begin // if (dataBuffer[WEIGHT_WIDTH] == 1'b1) 
                        case (dataBuffer01_re[SSAMPLE_WIDTH+WEIGHT_WIDTH -: SSAMPLE_WIDTH])
                            16'hFFFF: m01_axis_real_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= 16'hFFFF;
                            16'hEFFF: m01_axis_real_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= 16'hEFFF;
                            default:  m01_axis_real_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= dataBuffer01_re[SSAMPLE_WIDTH+WEIGHT_WIDTH -: SSAMPLE_WIDTH] + 1'b1;
                        endcase
                    end

                    dataBuffer01_im <= bw01_im*s01_axis_real_tdata[i*SSAMPLE_WIDTH +: SSAMPLE_WIDTH]
                        + bw01_re*s01_axis_imag_tdata[i*SSAMPLE_WIDTH +: SSAMPLE_WIDTH];
                    // rounding imaginary data using bit 8
                    if (dataBuffer01_im[WEIGHT_WIDTH] == 1'b0) begin
                        m01_axis_imag_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= dataBuffer01_im[SSAMPLE_WIDTH+WEIGHT_WIDTH -: SSAMPLE_WIDTH];
                    end
                    else begin // if (dataBuffer[WEIGHT_WIDTH] == 1'b1)
                        case (dataBuffer01_im[SSAMPLE_WIDTH+WEIGHT_WIDTH -: SSAMPLE_WIDTH])
                            16'hFFFF: m01_axis_imag_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= 16'hFFFF;
                            16'hEFFF: m01_axis_imag_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= 16'hEFFF;
                            default:  m01_axis_imag_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= dataBuffer01_im[SSAMPLE_WIDTH+WEIGHT_WIDTH -: SSAMPLE_WIDTH] + 1'b1;
                        endcase
                    end
                end
            end
            /*----------------------CHANNEL 01 NOT READY/VALID----------------------*/
            else begin 
                s01_axis_real_tready = 1'b0;       s01_axis_imag_tready = 1'b0;
                // invalid data, so output data is set to static value of 0
                m01_axis_real_s2mm_tdata <= 128'b0;
                m01_axis_imag_s2mm_tdata <= 128'b0;

                // output valid and output tkeep should be low
                m01_axis_real_s2mm_tvalid <= 1'b0; m01_axis_imag_s2mm_tvalid <= 1'b0;
                m01_axis_real_s2mm_tkeep <= 1'b0;  m01_axis_imag_s2mm_tkeep <= 1'b0;
            end
            /*------------------------CHANNEL 20 READY/VALID------------------------*/
            if (m20_axis_real_s2mm_tready && s20_axis_real_tvalid && m20_axis_imag_s2mm_tready && s20_axis_imag_tvalid) begin
                s20_axis_real_tready = 1'b1;       s20_axis_imag_tready = 1'b1;
                // tkeep and tvalid are now high (tkeep = 16'hffff, tvalid = 1'b1)
                m20_axis_real_s2mm_tkeep <= 16'hffff;   m20_axis_imag_s2mm_tkeep <= 16'hffff;
                m20_axis_real_s2mm_tvalid <= 1'b1;      m20_axis_imag_s2mm_tvalid <= 1'b1;

                // this for loop multiplies every eight bits by bWeights (it'll loop 16 times- 1 time per sample in tdata)
                for(i=0; i<samples; i = i+1) begin
                    // this can be a non-blocking assignment because there is a blocking assignment in the incrementing of i
                    // multiply by appropriate weight, accounting for complex/real parts of weight
                    dataBuffer20_re <= bw20_re*s20_axis_real_tdata[i*SSAMPLE_WIDTH +: SSAMPLE_WIDTH]
                        + bw20_im*s20_axis_imag_tdata[i*SSAMPLE_WIDTH +: SSAMPLE_WIDTH]; 
                    // rounding real data using bit 8
                    if (dataBuffer20_re[WEIGHT_WIDTH] == 1'b0) begin
                        m20_axis_real_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= dataBuffer20_re[SSAMPLE_WIDTH+WEIGHT_WIDTH -: SSAMPLE_WIDTH];
                    end
                    else begin // if (dataBuffer[WEIGHT_WIDTH] == 1'b1)
                        case (dataBuffer20_re[SSAMPLE_WIDTH+WEIGHT_WIDTH -: SSAMPLE_WIDTH])
                            16'hFFFF: m20_axis_real_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= 16'hFFFF;
                            16'hEFFF: m20_axis_real_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= 16'hEFFF;
                            default:  m20_axis_real_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= dataBuffer20_re[SSAMPLE_WIDTH+WEIGHT_WIDTH -: SSAMPLE_WIDTH] + 1'b1;
                        endcase
                    end

                    dataBuffer20_im <= bw20_im*s20_axis_real_tdata[i*SSAMPLE_WIDTH +: SSAMPLE_WIDTH]
                        + bw20_re*s20_axis_imag_tdata[i*SSAMPLE_WIDTH +: SSAMPLE_WIDTH];
                    // rounding imaginary data using bit 8
                    if (dataBuffer20_im[WEIGHT_WIDTH] == 1'b0) begin
                        m20_axis_imag_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= dataBuffer20_im[SSAMPLE_WIDTH+WEIGHT_WIDTH -: SSAMPLE_WIDTH];
                    end
                    else begin // if (dataBuffer[WEIGHT_WIDTH] == 1)
                        case (dataBuffer20_im[SSAMPLE_WIDTH+WEIGHT_WIDTH -: SSAMPLE_WIDTH])
                            16'hFFFF: m20_axis_imag_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= 16'hFFFF;
                            16'hEFFF: m20_axis_imag_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= 16'hEFFF;
                            default:  m20_axis_imag_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= dataBuffer20_im[SSAMPLE_WIDTH+WEIGHT_WIDTH -: SSAMPLE_WIDTH] + 1'b1;
                        endcase
                    end
                end
            end
            /*----------------------CHANNEL 20 NOT READY/VALID----------------------*/
            else begin 
                s20_axis_real_tready = 1'b0;       s20_axis_imag_tready = 1'b0;
                // invalid data, so output data is set to static value of 0
                m20_axis_real_s2mm_tdata <= 128'b0;
                m20_axis_imag_s2mm_tdata <= 128'b0;

                // output valid and output tkeep should be low
                m20_axis_real_s2mm_tvalid <= 1'b0; m20_axis_imag_s2mm_tvalid <= 1'b0;
                m20_axis_real_s2mm_tkeep <= 1'b0;  m20_axis_imag_s2mm_tkeep <= 1'b0;
            end
            /*------------------------CHANNEL 21 READY/VALID------------------------*/
            if (m21_axis_real_s2mm_tready && s21_axis_real_tvalid && m21_axis_imag_s2mm_tready && s21_axis_imag_tvalid) begin
                s21_axis_real_tready = 1'b1;       s21_axis_imag_tready = 1'b1;
                // tkeep and tvalid are now high (tkeep = 16'hffff, tvalid = 1'b1)
                m21_axis_real_s2mm_tkeep <= 16'hffff;   m21_axis_imag_s2mm_tkeep <= 16'hffff;
                m21_axis_real_s2mm_tvalid <= 1'b1;      m21_axis_imag_s2mm_tvalid <= 1'b1;

                // this for loop multiplies every eight bits by bWeights (it'll loop 16 times- 1 time per sample in tdata)
                for(i=0; i<samples; i = i+1) begin
                    // this can be a non-blocking assignment because there is a blocking assignment in the incrementing of i
                    // multiply by appropriate weight, accounting for complex/real parts of weight
                    dataBuffer21_re <= bw21_re*s21_axis_real_tdata[i*SSAMPLE_WIDTH +: SSAMPLE_WIDTH]
                        + bw21_im*s21_axis_imag_tdata[i*SSAMPLE_WIDTH +: SSAMPLE_WIDTH]; 
                    // rounding real data using bit 8
                    if (dataBuffer21_re[WEIGHT_WIDTH] == 1'b0) begin
                        m21_axis_real_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= dataBuffer21_re[SSAMPLE_WIDTH+WEIGHT_WIDTH -: SSAMPLE_WIDTH];
                    end
                    else begin // if (dataBuffer[WEIGHT_WIDTH] == 1'b1) 
                        case (dataBuffer21_re[SSAMPLE_WIDTH+WEIGHT_WIDTH -: SSAMPLE_WIDTH])
                            16'hFFFF: m21_axis_real_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= 16'hFFFF;
                            16'hEFFF: m21_axis_real_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= 16'hEFFF;
                            default:  m21_axis_real_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= dataBuffer21_re[SSAMPLE_WIDTH+WEIGHT_WIDTH -: SSAMPLE_WIDTH] + 1'b1;
                        endcase
                    end

                    dataBuffer21_im <= bw21_im*s21_axis_real_tdata[i*SSAMPLE_WIDTH +: SSAMPLE_WIDTH]
                        + bw21_re*s21_axis_imag_tdata[i*SSAMPLE_WIDTH +: SSAMPLE_WIDTH];
                    // rounding imaginary data using bit 8
                    if (dataBuffer21_im[WEIGHT_WIDTH] == 1'b0) begin
                        m21_axis_imag_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= dataBuffer21_im[SSAMPLE_WIDTH+WEIGHT_WIDTH -: SSAMPLE_WIDTH];
                    end
                    else begin // if (dataBuffer[WEIGHT_WIDTH] == 1'b1)
                        case (dataBuffer21_im[SSAMPLE_WIDTH+WEIGHT_WIDTH -: SSAMPLE_WIDTH])
                            16'hFFFF: m21_axis_imag_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= 16'hFFFF;
                            16'hEFFF: m21_axis_imag_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= 16'hEFFF;
                            default:  m21_axis_imag_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= dataBuffer21_im[SSAMPLE_WIDTH+WEIGHT_WIDTH -: SSAMPLE_WIDTH] + 1'b1;
                        endcase
                    end
                end
            end
            /*----------------------CHANNEL 21 NOT READY/VALID----------------------*/
            else begin 
                s21_axis_real_tready = 1'b0;       s21_axis_imag_tready = 1'b0;
                // invalid data, so output data is set to static value of 0
                m21_axis_real_s2mm_tdata <= 128'b0;
                m21_axis_imag_s2mm_tdata <= 128'b0;

                // output valid and output tkeep should be low
                m21_axis_real_s2mm_tvalid <= 1'b0; m21_axis_imag_s2mm_tvalid <= 1'b0;
                m21_axis_real_s2mm_tkeep <= 1'b0;  m21_axis_imag_s2mm_tkeep <= 1'b0;
            end

            /* 1. This implementation of the Adder assumes that if one channel has valid data, so do the rest of the channels
             * The data it produces should be accurate, but given how I'm rounding the data, the firmware may be faster
             * and more precise if I only sum the data if two or more channels have valid data.
             *
             * 2. Additionally, the data may be more precise if I round based on how many channels have valid data (that we are summing)
             */
            if((s00_axis_real_tready && s00_axis_imag_tready) || (s01_axis_real_tready && s01_axis_imag_tready)  ||
               (s20_axis_real_tready && s20_axis_imag_tready) || (s21_axis_real_tready && s21_axis_imag_tready)) begin
                // this for loop multiplies every eight bits by bWeights (it'll loop 16 times- 1 time per sample in tdata)
                for(i=0; i<samples; i = i+1) begin
                    // this can be a non-blocking assignment because there is a blocking assignment in the incrementing of i
                    dataBuffer_SumRe <= m00_axis_real_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] + m01_axis_real_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH]
                        + m20_axis_real_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] + m21_axis_real_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH];
                    if (dataBuffer_SumRe[2] == 1'b1) begin // round up
                        case (dataBuffer_SumRe[MSAMPLE_WIDTH+2 -: MSAMPLE_WIDTH])
                            16'hFFFF: m00_axis_real_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= 16'hFFFF;
                            16'hEFFF: m00_axis_real_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= 16'hEFFF;
                            default:  m00_axis_real_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= dataBuffer_SumRe[MSAMPLE_WIDTH+2 -: MSAMPLE_WIDTH] + 1'b1;
                        endcase
                    end
                    else begin // round down
                        m00_axis_real_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= dataBuffer_SumRe[MSAMPLE_WIDTH+2 -: MSAMPLE_WIDTH];
                    end

                    dataBuffer_SumIm <= m00_axis_imag_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] + m01_axis_imag_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH]
                        + m20_axis_imag_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] + m21_axis_imag_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH];
                    if (dataBuffer_SumIm[2] == 1'b1) begin // round up
                        case (dataBuffer_SumIm[MSAMPLE_WIDTH+2 -: MSAMPLE_WIDTH])
                            16'hFFFF: m00_axis_imag_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= 16'hFFFF;
                            16'hEFFF: m00_axis_imag_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= 16'hEFFF;
                            default:  m00_axis_imag_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= dataBuffer_SumIm[MSAMPLE_WIDTH+2 -: MSAMPLE_WIDTH] + 1'b1;
                        endcase
                    end
                    else begin // round down
                        m00_axis_imag_s2mm_tdata[i*MSAMPLE_WIDTH +: MSAMPLE_WIDTH] <= dataBuffer_SumIm[MSAMPLE_WIDTH+2 -: MSAMPLE_WIDTH];
                    end
                end
            end
         end
    end
endmodule
