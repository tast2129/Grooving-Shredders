hsfgdg
